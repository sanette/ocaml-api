../search_icon.sv